-----------------------------------------------------------------------
-- Project: CiM-Tile HW Design/implementation                        --
-- File	  : instruction_memory_1.vhd                                 --
-- Author : Remon van Duijnen (R.F.J.vanDuijnen@student.tudelft.nl)  --
-- Version: 1.0														 --
-----------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.math_real.all;
use ieee.numeric_std.all;

entity instruction_memory_1 is
	generic(inst_size : integer;
			PC_size   : integer;
			mem_size  : integer);
	port( i_PC : in std_logic_vector(PC_size - 1 downto 0);

		  o_inst : out std_logic_vector(inst_size * 8 - 1 downto 0)
);
end instruction_memory_1;

architecture behavioural of instruction_memory_1 is

	type inst_array_type is array (inst_size - 1 downto 0) of std_logic_vector(7 downto 0);
	type mem_array_type is array (mem_size - 1 downto 0) of std_logic_vector(7 downto 0);
	signal inst_array : inst_array_type;
	
	-- This constant should contain the stage 1 instruction bytes generated by the inst2HDL script (from compiler project)
	constant instruction_mem : mem_array_type := (

	0 => "01000000",
	1 => "00000000",
	2 => "01010000",
	3 => "00000000",
	4 => "11010000",
	5 => "00010000",
	6 => "00000000",
	7 => "00000001",
	8 => "01100000",
	9 => "00000011",
	10 => "01100000",
	11 => "00000010",
	12 => "01100000",
	13 => "00000001",
	14 => "01100000",
	15 => "00000000",
	16 => "10100000",
	17 => "10000000",
	18 => "01010000",
	19 => "00000000",
	20 => "11010000",
	21 => "00010000",
	22 => "00000000",
	23 => "00000010",
	24 => "01100000",
	25 => "00000011",
	26 => "01100000",
	27 => "00000010",
	28 => "01100000",
	29 => "00000001",
	30 => "01100000",
	31 => "00000000",
	32 => "10100000",
	33 => "10000000",
	34 => "01010000",
	35 => "00000000",
	36 => "11010000",
	37 => "00010000",
	38 => "00000000",
	39 => "00000100",
	40 => "01100000",
	41 => "00000011",
	42 => "01100000",
	43 => "00000010",
	44 => "01100000",
	45 => "00000001",
	46 => "01100000",
	47 => "00000000",
	48 => "10100000",
	49 => "10000000",
	50 => "01010000",
	51 => "00000000",
	52 => "11010000",
	53 => "00010000",
	54 => "00000000",
	55 => "00001000",
	56 => "01100000",
	57 => "00000011",
	58 => "01100000",
	59 => "00000010",
	60 => "01100000",
	61 => "00000001",
	62 => "01100000",
	63 => "00000000",
	64 => "10100000",
	65 => "10000000",
	66 => "01010000",
	67 => "00000000",
	68 => "11010000",
	69 => "00010000",
	70 => "00000000",
	71 => "00010000",
	72 => "01100000",
	73 => "00000011",
	74 => "01100000",
	75 => "00000010",
	76 => "01100000",
	77 => "00000001",
	78 => "01100000",
	79 => "00000000",
	80 => "10100000",
	81 => "10000000",
	82 => "01010000",
	83 => "00000000",
	84 => "11010000",
	85 => "00010000",
	86 => "00000000",
	87 => "00100000",
	88 => "01100000",
	89 => "00000011",
	90 => "01100000",
	91 => "00000010",
	92 => "01100000",
	93 => "00000001",
	94 => "01100000",
	95 => "00000000",
	96 => "10100000",
	97 => "10000000",
	98 => "01010000",
	99 => "00000000",
	100 => "11010000",
	101 => "00010000",
	102 => "00000000",
	103 => "01000000",
	104 => "01100000",
	105 => "00000011",
	106 => "01100000",
	107 => "00000010",
	108 => "01100000",
	109 => "00000001",
	110 => "01100000",
	111 => "00000000",
	112 => "10100000",
	113 => "10000000",
	114 => "01010000",
	115 => "00000000",
	116 => "11010000",
	117 => "00010000",
	118 => "00000000",
	119 => "10000000",
	120 => "01100000",
	121 => "00000011",
	122 => "01100000",
	123 => "00000010",
	124 => "01100000",
	125 => "00000001",
	126 => "01100000",
	127 => "00000000",
	128 => "10100000",
	129 => "10000000",
	130 => "01010000",
	131 => "00000000",
	132 => "11010000",
	133 => "00010000",
	134 => "00000001",
	135 => "00000001",
	136 => "01100000",
	137 => "00000011",
	138 => "01100000",
	139 => "00000010",
	140 => "01100000",
	141 => "00000001",
	142 => "01100000",
	143 => "00000000",
	144 => "10100000",
	145 => "10000000",
	146 => "01010000",
	147 => "00000000",
	148 => "11010000",
	149 => "00010000",
	150 => "00000001",
	151 => "00000010",
	152 => "01100000",
	153 => "00000011",
	154 => "01100000",
	155 => "00000010",
	156 => "01100000",
	157 => "00000001",
	158 => "01100000",
	159 => "00000000",
	160 => "10100000",
	161 => "10000000",
	162 => "01010000",
	163 => "00000000",
	164 => "11010000",
	165 => "00010000",
	166 => "00000001",
	167 => "00000100",
	168 => "01100000",
	169 => "00000011",
	170 => "01100000",
	171 => "00000010",
	172 => "01100000",
	173 => "00000001",
	174 => "01100000",
	175 => "00000000",
	176 => "10100000",
	177 => "10000000",
	178 => "01010000",
	179 => "00000000",
	180 => "11010000",
	181 => "00010000",
	182 => "00000001",
	183 => "00001000",
	184 => "01100000",
	185 => "00000011",
	186 => "01100000",
	187 => "00000010",
	188 => "01100000",
	189 => "00000001",
	190 => "01100000",
	191 => "00000000",
	192 => "10100000",
	193 => "10000000",
	194 => "01010000",
	195 => "00000000",
	196 => "11010000",
	197 => "00010000",
	198 => "00000001",
	199 => "00010000",
	200 => "01100000",
	201 => "00000011",
	202 => "01100000",
	203 => "00000010",
	204 => "01100000",
	205 => "00000001",
	206 => "01100000",
	207 => "00000000",
	208 => "10100000",
	209 => "10000000",
	210 => "01010000",
	211 => "00000000",
	212 => "11010000",
	213 => "00010000",
	214 => "00000001",
	215 => "00100000",
	216 => "01100000",
	217 => "00000011",
	218 => "01100000",
	219 => "00000010",
	220 => "01100000",
	221 => "00000001",
	222 => "01100000",
	223 => "00000000",
	224 => "10100000",
	225 => "10000000",
	226 => "01010000",
	227 => "00000000",
	228 => "11010000",
	229 => "00010000",
	230 => "00000001",
	231 => "01000000",
	232 => "01100000",
	233 => "00000011",
	234 => "01100000",
	235 => "00000010",
	236 => "01100000",
	237 => "00000001",
	238 => "01100000",
	239 => "00000000",
	240 => "10100000",
	241 => "10000000",
	242 => "01010000",
	243 => "00000000",
	244 => "11010000",
	245 => "00010000",
	246 => "00000001",
	247 => "10000000",
	248 => "01100000",
	249 => "00000011",
	250 => "01100000",
	251 => "00000010",
	252 => "01100000",
	253 => "00000001",
	254 => "01100000",
	255 => "00000000",
	256 => "10100000",
	257 => "10000000",
	258 => "01010000",
	259 => "00000000",
	260 => "11010000",
	261 => "00010000",
	262 => "00000010",
	263 => "00000001",
	264 => "01100000",
	265 => "00000011",
	266 => "01100000",
	267 => "00000010",
	268 => "01100000",
	269 => "00000001",
	270 => "01100000",
	271 => "00000000",
	272 => "10100000",
	273 => "10000000",
	274 => "01010000",
	275 => "00000000",
	276 => "11010000",
	277 => "00010000",
	278 => "00000010",
	279 => "00000010",
	280 => "01100000",
	281 => "00000011",
	282 => "01100000",
	283 => "00000010",
	284 => "01100000",
	285 => "00000001",
	286 => "01100000",
	287 => "00000000",
	288 => "10100000",
	289 => "10000000",
	290 => "01010000",
	291 => "00000000",
	292 => "11010000",
	293 => "00010000",
	294 => "00000010",
	295 => "00000100",
	296 => "01100000",
	297 => "00000011",
	298 => "01100000",
	299 => "00000010",
	300 => "01100000",
	301 => "00000001",
	302 => "01100000",
	303 => "00000000",
	304 => "10100000",
	305 => "10000000",
	306 => "01010000",
	307 => "00000000",
	308 => "11010000",
	309 => "00010000",
	310 => "00000010",
	311 => "00001000",
	312 => "01100000",
	313 => "00000011",
	314 => "01100000",
	315 => "00000010",
	316 => "01100000",
	317 => "00000001",
	318 => "01100000",
	319 => "00000000",
	320 => "10100000",
	321 => "10000000",
	322 => "01010000",
	323 => "00000000",
	324 => "11010000",
	325 => "00010000",
	326 => "00000010",
	327 => "00010000",
	328 => "01100000",
	329 => "00000011",
	330 => "01100000",
	331 => "00000010",
	332 => "01100000",
	333 => "00000001",
	334 => "01100000",
	335 => "00000000",
	336 => "10100000",
	337 => "10000000",
	338 => "01010000",
	339 => "00000000",
	340 => "11010000",
	341 => "00010000",
	342 => "00000010",
	343 => "00100000",
	344 => "01100000",
	345 => "00000011",
	346 => "01100000",
	347 => "00000010",
	348 => "01100000",
	349 => "00000001",
	350 => "01100000",
	351 => "00000000",
	352 => "10100000",
	353 => "10000000",
	354 => "01010000",
	355 => "00000000",
	356 => "11010000",
	357 => "00010000",
	358 => "00000010",
	359 => "01000000",
	360 => "01100000",
	361 => "00000011",
	362 => "01100000",
	363 => "00000010",
	364 => "01100000",
	365 => "00000001",
	366 => "01100000",
	367 => "00000000",
	368 => "10100000",
	369 => "10000000",
	370 => "01010000",
	371 => "00000000",
	372 => "11010000",
	373 => "00010000",
	374 => "00000010",
	375 => "10000000",
	376 => "01100000",
	377 => "00000011",
	378 => "01100000",
	379 => "00000010",
	380 => "01100000",
	381 => "00000001",
	382 => "01100000",
	383 => "00000000",
	384 => "10100000",
	385 => "10000000",
	386 => "01010000",
	387 => "00000000",
	388 => "11010000",
	389 => "00010000",
	390 => "00000011",
	391 => "00000001",
	392 => "01100000",
	393 => "00000011",
	394 => "01100000",
	395 => "00000010",
	396 => "01100000",
	397 => "00000001",
	398 => "01100000",
	399 => "00000000",
	400 => "10100000",
	401 => "10000000",
	402 => "01010000",
	403 => "00000000",
	404 => "11010000",
	405 => "00010000",
	406 => "00000011",
	407 => "00000010",
	408 => "01100000",
	409 => "00000011",
	410 => "01100000",
	411 => "00000010",
	412 => "01100000",
	413 => "00000001",
	414 => "01100000",
	415 => "00000000",
	416 => "10100000",
	417 => "10000000",
	418 => "01010000",
	419 => "00000000",
	420 => "11010000",
	421 => "00010000",
	422 => "00000011",
	423 => "00000100",
	424 => "01100000",
	425 => "00000011",
	426 => "01100000",
	427 => "00000010",
	428 => "01100000",
	429 => "00000001",
	430 => "01100000",
	431 => "00000000",
	432 => "10100000",
	433 => "10000000",
	434 => "01010000",
	435 => "00000000",
	436 => "11010000",
	437 => "00010000",
	438 => "00000011",
	439 => "00001000",
	440 => "01100000",
	441 => "00000011",
	442 => "01100000",
	443 => "00000010",
	444 => "01100000",
	445 => "00000001",
	446 => "01100000",
	447 => "00000000",
	448 => "10100000",
	449 => "10000000",
	450 => "01010000",
	451 => "00000000",
	452 => "11010000",
	453 => "00010000",
	454 => "00000011",
	455 => "00010000",
	456 => "01100000",
	457 => "00000011",
	458 => "01100000",
	459 => "00000010",
	460 => "01100000",
	461 => "00000001",
	462 => "01100000",
	463 => "00000000",
	464 => "10100000",
	465 => "10000000",
	466 => "01010000",
	467 => "00000000",
	468 => "11010000",
	469 => "00010000",
	470 => "00000011",
	471 => "00100000",
	472 => "01100000",
	473 => "00000011",
	474 => "01100000",
	475 => "00000010",
	476 => "01100000",
	477 => "00000001",
	478 => "01100000",
	479 => "00000000",
	480 => "10100000",
	481 => "10000000",
	482 => "01010000",
	483 => "00000000",
	484 => "11010000",
	485 => "00010000",
	486 => "00000011",
	487 => "01000000",
	488 => "01100000",
	489 => "00000011",
	490 => "01100000",
	491 => "00000010",
	492 => "01100000",
	493 => "00000001",
	494 => "01100000",
	495 => "00000000",
	496 => "10100000",
	497 => "10000000",
	498 => "01010000",
	499 => "00000000",
	500 => "11010000",
	501 => "00010000",
	502 => "00000011",
	503 => "10000000",
	504 => "01100000",
	505 => "00000011",
	506 => "01100000",
	507 => "00000010",
	508 => "01100000",
	509 => "00000001",
	510 => "01100000",
	511 => "00000000",
	512 => "10100000",
	513 => "10000000",
	514 => "01010000",
	515 => "00000111",
	516 => "11100000",
	517 => "11000000",
	518 => "10000000",
	519 => "10010000",
	520 => "01010000",
	521 => "00000111",
	522 => "11100000",
	523 => "10000000",
	524 => "10010000",
	525 => "01010000",
	526 => "00000111",
	527 => "11100000",
	528 => "10000000",
	529 => "10010000",
	530 => "01010000",
	531 => "00000111",
	532 => "11100000",
	533 => "10000000",
	534 => "10010000",
	535 => "01010000",
	536 => "00000111",
	537 => "11100000",
	538 => "10000000",
	539 => "10010000",
	540 => "01010000",
	541 => "00000111",
	542 => "11100000",
	543 => "10000000",
	544 => "10010000",
	545 => "01010000",
	546 => "00000111",
	547 => "11100000",
	548 => "10000000",
	549 => "10010000",
	550 => "01010000",
	551 => "00000111",
	552 => "11100000",
	553 => "10000000",
	554 => "10010000",
	555 => "01010000",
	556 => "00000111",
	557 => "11100000",
	558 => "10000000",
	559 => "10010000",
	560 => "01010000",
	561 => "00000111",
	562 => "11100000",
	563 => "10000000",
	564 => "10010000",
	565 => "01010000",
	566 => "00000111",
	567 => "11100000",
	568 => "10000000",
	569 => "10010000",
	570 => "01010000",
	571 => "00000111",
	572 => "11100000",
	573 => "10000000",
	574 => "10010000",
	575 => "01010000",
	576 => "00000111",
	577 => "11100000",
	578 => "10000000",
	579 => "10010000",
	580 => "01010000",
	581 => "00000111",
	582 => "11100000",
	583 => "10000000",
	584 => "10010000",
	585 => "01010000",
	586 => "00000111",
	587 => "11100000",
	588 => "10000000",
	589 => "10010000",
	590 => "01010000",
	591 => "00000111",
	592 => "11100000",
	593 => "10000000",
	594 => "10010000",
	595 => "01010000",
	596 => "00000111",
	597 => "11100000",
	598 => "10000000",
	599 => "10010000",
	600 => "01010000",
	601 => "00000111",
	602 => "11100000",
	603 => "10000000",
	604 => "10010000",
	605 => "01010000",
	606 => "00000111",
	607 => "11100000",
	608 => "10000000",
	609 => "10010000",
	610 => "01010000",
	611 => "00000111",
	612 => "11100000",
	613 => "10000000",
	614 => "10010000",
	615 => "01010000",
	616 => "00000111",
	617 => "11100000",
	618 => "10000000",
	619 => "10010000",
	620 => "01010000",
	621 => "00000111",
	622 => "11100000",
	623 => "10000000",
	624 => "10010000",
	625 => "01010000",
	626 => "00000111",
	627 => "11100000",
	628 => "10000000",
	629 => "10010000",
	630 => "01010000",
	631 => "00000111",
	632 => "11100000",
	633 => "10000000",
	634 => "10010000",
	635 => "01010000",
	636 => "00000111",
	637 => "11100000",
	638 => "10000000",
	639 => "10010000",
	640 => "01010000",
	641 => "00000111",
	642 => "11100000",
	643 => "10000000",
	644 => "10010000",
	645 => "01010000",
	646 => "00000111",
	647 => "11100000",
	648 => "10000000",
	649 => "10010000",
	650 => "01010000",
	651 => "00000111",
	652 => "11100000",
	653 => "10000000",
	654 => "10010000",
	655 => "01010000",
	656 => "00000111",
	657 => "11100000",
	658 => "10000000",
	659 => "10010000",
	660 => "01010000",
	661 => "00000111",
	662 => "11100000",
	663 => "10000000",
	664 => "10010000",
	665 => "01010000",
	666 => "00000111",
	667 => "11100000",
	668 => "10000000",
	669 => "10010000",
	670 => "01010000",
	671 => "00000111",
	672 => "11100000",
	673 => "10000000",
	674 => "10010000",
	675 => "00000000",
	others => "00000000"

);

begin

    -- fetch instruction based on PC
	process(i_PC)
	begin
		for i in inst_size - 1 downto 0 loop
			inst_array(inst_size - (i+1))	<= instruction_mem(to_integer(unsigned(i_PC))+i);
		end loop;

	end process;

    -- put instruction into array of bytes
G0: for i in inst_size - 1 downto 0 generate
G1: 	for j in 7 downto 0 generate
			o_inst(i * 8 + j) <= inst_array(i)(j);
		end generate;
	end generate;
	
 end behavioural;