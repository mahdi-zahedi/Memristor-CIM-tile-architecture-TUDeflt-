-----------------------------------------------------------------------
-- Project: CiM-Tile HW Design/implementation                        --
-- File	  : instruction_memory_2.vhd                                 --
-- Author : Remon van Duijnen (R.F.J.vanDuijnen@student.tudelft.nl)  --
-- Version: 1.0														 --
-----------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.math_real.all;
use ieee.numeric_std.all;

entity instruction_memory_2 is
	generic(inst_size : integer;
			PC_size   : integer;
			mem_size  : integer);
	port( i_PC : in std_logic_vector(PC_size - 1 downto 0);

		  o_inst : out std_logic_vector(inst_size * 8 - 1 downto 0)
);
end instruction_memory_2;

architecture behavioural of instruction_memory_2 is

	type inst_array_type is array (inst_size - 1 downto 0) of std_logic_vector(7 downto 0);
	type mem_array_type is array (mem_size - 1 downto 0) of std_logic_vector(7 downto 0);

	signal inst_array : inst_array_type;
	
	-- This constant should contain the stage 2 instruction bytes generated by the inst2HDL script (from compiler project)
	constant  instruction_mem : mem_array_type := (

	0 => "11000000",
	1 => "00010000",
	2 => "11000000",
	3 => "00000000",
	4 => "00010000",
	5 => "11000000",
	6 => "00000001",
	7 => "00010000",
	8 => "11000000",
	9 => "00000010",
	10 => "00010000",
	11 => "11000000",
	12 => "00000011",
	13 => "00010000",
	14 => "11000000",
	15 => "00000100",
	16 => "00010000",
	17 => "11000000",
	18 => "00000101",
	19 => "00010000",
	20 => "11000000",
	21 => "00000110",
	22 => "00010000",
	23 => "11000000",
	24 => "00000111",
	25 => "10000000",
	26 => "11010000",
	27 => "11000000",
	28 => "01000000",
	29 => "00000000",
	30 => "00000001",
	31 => "11010000",
	32 => "11000000",
	33 => "01000000",
	34 => "00000000",
	35 => "00000001",
	36 => "11010000",
	37 => "11000000",
	38 => "01000000",
	39 => "00000000",
	40 => "00000001",
	41 => "11010000",
	42 => "11000000",
	43 => "01000000",
	44 => "00000000",
	45 => "00000001",
	46 => "11010000",
	47 => "11000000",
	48 => "01000000",
	49 => "00000000",
	50 => "00000001",
	51 => "11010000",
	52 => "11000000",
	53 => "01000000",
	54 => "00000000",
	55 => "00000001",
	56 => "11010000",
	57 => "11000000",
	58 => "01000000",
	59 => "00000000",
	60 => "00000001",
	61 => "11010000",
	62 => "11100000",
	63 => "11000000",
	64 => "00010000",
	65 => "11000000",
	66 => "00001000",
	67 => "00010000",
	68 => "11000000",
	69 => "00001001",
	70 => "00010000",
	71 => "11000000",
	72 => "00001010",
	73 => "00010000",
	74 => "11000000",
	75 => "00001011",
	76 => "00010000",
	77 => "11000000",
	78 => "00001100",
	79 => "00010000",
	80 => "11000000",
	81 => "00001101",
	82 => "00010000",
	83 => "11000000",
	84 => "00001110",
	85 => "00010000",
	86 => "11000000",
	87 => "00001111",
	88 => "10000000",
	89 => "11010000",
	90 => "11000000",
	91 => "01000000",
	92 => "00000000",
	93 => "01000000",
	94 => "11010000",
	95 => "11000000",
	96 => "01000000",
	97 => "00000000",
	98 => "01000000",
	99 => "11010000",
	100 => "11000000",
	101 => "01000000",
	102 => "00000000",
	103 => "01000000",
	104 => "11010000",
	105 => "11000000",
	106 => "01000000",
	107 => "00000000",
	108 => "01000000",
	109 => "11010000",
	110 => "11000000",
	111 => "01000000",
	112 => "00000000",
	113 => "01000000",
	114 => "11010000",
	115 => "11000000",
	116 => "01000000",
	117 => "00000000",
	118 => "01000000",
	119 => "11010000",
	120 => "11000000",
	121 => "01000000",
	122 => "00000000",
	123 => "01000000",
	124 => "11010000",
	125 => "11100000",
	126 => "11000000",
	127 => "00010000",
	128 => "11000000",
	129 => "00000000",
	130 => "00010000",
	131 => "11000000",
	132 => "00000001",
	133 => "00010000",
	134 => "11000000",
	135 => "00000010",
	136 => "00010000",
	137 => "11000000",
	138 => "00000011",
	139 => "00010000",
	140 => "11000000",
	141 => "00000100",
	142 => "00010000",
	143 => "11000000",
	144 => "00000101",
	145 => "00010000",
	146 => "11000000",
	147 => "00000110",
	148 => "00010000",
	149 => "11000000",
	150 => "00000111",
	151 => "10000000",
	152 => "11010000",
	153 => "11000000",
	154 => "01000000",
	155 => "00000000",
	156 => "01111111",
	157 => "11010000",
	158 => "11000000",
	159 => "01000000",
	160 => "00000000",
	161 => "01111111",
	162 => "11010000",
	163 => "11000000",
	164 => "01000000",
	165 => "00000000",
	166 => "01111111",
	167 => "11010000",
	168 => "11000000",
	169 => "01000000",
	170 => "00000000",
	171 => "01111111",
	172 => "11010000",
	173 => "11000000",
	174 => "01000000",
	175 => "00000000",
	176 => "01111111",
	177 => "11010000",
	178 => "11000000",
	179 => "01000000",
	180 => "00000000",
	181 => "01111111",
	182 => "11010000",
	183 => "11000000",
	184 => "01000000",
	185 => "00000000",
	186 => "01111111",
	187 => "11010000",
	188 => "11100000",
	189 => "11000000",
	190 => "00010000",
	191 => "11000000",
	192 => "00001000",
	193 => "00010000",
	194 => "11000000",
	195 => "00001001",
	196 => "00010000",
	197 => "11000000",
	198 => "00001010",
	199 => "00010000",
	200 => "11000000",
	201 => "00001011",
	202 => "00010000",
	203 => "11000000",
	204 => "00001100",
	205 => "00010000",
	206 => "11000000",
	207 => "00001101",
	208 => "00010000",
	209 => "11000000",
	210 => "00001110",
	211 => "00010000",
	212 => "11000000",
	213 => "00001111",
	214 => "10000000",
	215 => "11010000",
	216 => "11000000",
	217 => "01000000",
	218 => "00000000",
	219 => "10111110",
	220 => "11010000",
	221 => "11000000",
	222 => "01000000",
	223 => "00000000",
	224 => "10111110",
	225 => "11010000",
	226 => "11000000",
	227 => "01000000",
	228 => "00000000",
	229 => "10111110",
	230 => "11010000",
	231 => "11000000",
	232 => "01000000",
	233 => "00000000",
	234 => "10111110",
	235 => "11010000",
	236 => "11000000",
	237 => "01000000",
	238 => "00000000",
	239 => "10111110",
	240 => "11010000",
	241 => "11000000",
	242 => "01000000",
	243 => "00000000",
	244 => "10111110",
	245 => "11010000",
	246 => "11000000",
	247 => "01000000",
	248 => "00000000",
	249 => "10111110",
	250 => "11010000",
	251 => "11100000",
	252 => "00000000",
	others => "00000000"

);

begin

    -- fetch next instruction based on PC
	process(i_PC)
	begin
		for i in inst_size - 1 downto 0 loop
			inst_array(inst_size - (i + 1))	<= instruction_mem(to_integer(unsigned(i_PC))+i);
		end loop;
	end process;

    -- put the instruction into an array of bytes
G0: for i in inst_size - 1 downto 0 generate
G1: 	for j in 7 downto 0 generate
			o_inst(i * 8 + j) <= inst_array(i)(j);
		end generate;
	end generate;
	


end behavioural;